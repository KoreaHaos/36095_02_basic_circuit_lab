** Profile: "SCHEMATIC1-lab2part2sim1"  [ C:\Users\Ben-Setup\Desktop\test\1\week2_lab-PSpiceFiles\SCHEMATIC1\lab2part2sim1.sim ] 

** Creating circuit file "lab2part2sim1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Ben-Setup\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V2 0V 1V 0.1V 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
