** Profile: "SCHEMATIC1-lab1part1sim1"  [ C:\Users\Ben-Setup\Desktop\test_workspace\lab1part1-PSpiceFiles\SCHEMATIC1\lab1part1sim1.sim ] 

** Creating circuit file "lab1part1sim1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Ben-Setup\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V1 0V 6V .1V 
+ LIN I_I1 0 5mA 0.5mA 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
